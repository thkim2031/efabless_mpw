VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLA_16
  CLASS BLOCK ;
  FOREIGN CLA_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 79.165 BY 89.885 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END CIN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END CLK
  PIN COUT_FINAL
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END COUT_FINAL
  PIN OPA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END OPA[0]
  PIN OPA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 85.885 0.370 89.885 ;
    END
  END OPA[10]
  PIN OPA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 37.440 79.165 38.040 ;
    END
  END OPA[11]
  PIN OPA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 85.885 64.770 89.885 ;
    END
  END OPA[12]
  PIN OPA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END OPA[13]
  PIN OPA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 10.240 79.165 10.840 ;
    END
  END OPA[14]
  PIN OPA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 85.885 51.890 89.885 ;
    END
  END OPA[15]
  PIN OPA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 3.440 79.165 4.040 ;
    END
  END OPA[1]
  PIN OPA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END OPA[2]
  PIN OPA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 17.040 79.165 17.640 ;
    END
  END OPA[3]
  PIN OPA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 85.885 6.810 89.885 ;
    END
  END OPA[4]
  PIN OPA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 23.840 79.165 24.440 ;
    END
  END OPA[5]
  PIN OPA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END OPA[6]
  PIN OPA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 85.885 32.570 89.885 ;
    END
  END OPA[7]
  PIN OPA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END OPA[8]
  PIN OPA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END OPA[9]
  PIN OPB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END OPB[0]
  PIN OPB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END OPB[10]
  PIN OPB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END OPB[11]
  PIN OPB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 64.640 79.165 65.240 ;
    END
  END OPB[12]
  PIN OPB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END OPB[13]
  PIN OPB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 85.885 45.450 89.885 ;
    END
  END OPB[14]
  PIN OPB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 85.885 26.130 89.885 ;
    END
  END OPB[15]
  PIN OPB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 85.040 79.165 85.640 ;
    END
  END OPB[1]
  PIN OPB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 71.440 79.165 72.040 ;
    END
  END OPB[2]
  PIN OPB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 51.040 79.165 51.640 ;
    END
  END OPB[3]
  PIN OPB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 85.885 58.330 89.885 ;
    END
  END OPB[4]
  PIN OPB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END OPB[5]
  PIN OPB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END OPB[6]
  PIN OPB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END OPB[7]
  PIN OPB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 78.240 79.165 78.840 ;
    END
  END OPB[8]
  PIN OPB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END OPB[9]
  PIN PHI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 57.840 79.165 58.440 ;
    END
  END PHI
  PIN SUM_FINAL[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END SUM_FINAL[0]
  PIN SUM_FINAL[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 85.885 39.010 89.885 ;
    END
  END SUM_FINAL[10]
  PIN SUM_FINAL[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 30.640 79.165 31.240 ;
    END
  END SUM_FINAL[11]
  PIN SUM_FINAL[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END SUM_FINAL[12]
  PIN SUM_FINAL[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END SUM_FINAL[13]
  PIN SUM_FINAL[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END SUM_FINAL[14]
  PIN SUM_FINAL[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END SUM_FINAL[15]
  PIN SUM_FINAL[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END SUM_FINAL[1]
  PIN SUM_FINAL[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 85.885 77.650 89.885 ;
    END
  END SUM_FINAL[2]
  PIN SUM_FINAL[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 85.885 71.210 89.885 ;
    END
  END SUM_FINAL[3]
  PIN SUM_FINAL[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 85.885 13.250 89.885 ;
    END
  END SUM_FINAL[4]
  PIN SUM_FINAL[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 85.885 19.690 89.885 ;
    END
  END SUM_FINAL[5]
  PIN SUM_FINAL[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END SUM_FINAL[6]
  PIN SUM_FINAL[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END SUM_FINAL[7]
  PIN SUM_FINAL[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END SUM_FINAL[8]
  PIN SUM_FINAL[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 75.165 44.240 79.165 44.840 ;
    END
  END SUM_FINAL[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 21.740 10.640 23.340 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.760 10.640 40.360 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 55.780 10.640 57.380 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.800 10.640 74.400 79.120 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 13.230 10.640 14.830 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 30.250 10.640 31.850 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 47.270 10.640 48.870 79.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.290 10.640 65.890 79.120 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 73.600 78.965 ;
      LAYER met1 ;
        RECT 0.070 5.480 77.670 79.120 ;
      LAYER met2 ;
        RECT 0.650 85.605 6.250 85.885 ;
        RECT 7.090 85.605 12.690 85.885 ;
        RECT 13.530 85.605 19.130 85.885 ;
        RECT 19.970 85.605 25.570 85.885 ;
        RECT 26.410 85.605 32.010 85.885 ;
        RECT 32.850 85.605 38.450 85.885 ;
        RECT 39.290 85.605 44.890 85.885 ;
        RECT 45.730 85.605 51.330 85.885 ;
        RECT 52.170 85.605 57.770 85.885 ;
        RECT 58.610 85.605 64.210 85.885 ;
        RECT 65.050 85.605 70.650 85.885 ;
        RECT 71.490 85.605 77.090 85.885 ;
        RECT 0.100 4.280 77.640 85.605 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 19.130 4.280 ;
        RECT 19.970 3.555 25.570 4.280 ;
        RECT 26.410 3.555 32.010 4.280 ;
        RECT 32.850 3.555 38.450 4.280 ;
        RECT 39.290 3.555 44.890 4.280 ;
        RECT 45.730 3.555 51.330 4.280 ;
        RECT 52.170 3.555 57.770 4.280 ;
        RECT 58.610 3.555 64.210 4.280 ;
        RECT 65.050 3.555 70.650 4.280 ;
        RECT 71.490 3.555 77.090 4.280 ;
      LAYER met3 ;
        RECT 4.400 84.640 74.765 85.505 ;
        RECT 4.000 79.240 76.050 84.640 ;
        RECT 4.400 77.840 74.765 79.240 ;
        RECT 4.000 72.440 76.050 77.840 ;
        RECT 4.400 71.040 74.765 72.440 ;
        RECT 4.000 65.640 76.050 71.040 ;
        RECT 4.400 64.240 74.765 65.640 ;
        RECT 4.000 58.840 76.050 64.240 ;
        RECT 4.400 57.440 74.765 58.840 ;
        RECT 4.000 52.040 76.050 57.440 ;
        RECT 4.400 50.640 74.765 52.040 ;
        RECT 4.000 45.240 76.050 50.640 ;
        RECT 4.400 43.840 74.765 45.240 ;
        RECT 4.000 38.440 76.050 43.840 ;
        RECT 4.400 37.040 74.765 38.440 ;
        RECT 4.000 31.640 76.050 37.040 ;
        RECT 4.400 30.240 74.765 31.640 ;
        RECT 4.000 24.840 76.050 30.240 ;
        RECT 4.400 23.440 74.765 24.840 ;
        RECT 4.000 18.040 76.050 23.440 ;
        RECT 4.400 16.640 74.765 18.040 ;
        RECT 4.000 11.240 76.050 16.640 ;
        RECT 4.400 9.840 74.765 11.240 ;
        RECT 4.000 4.440 76.050 9.840 ;
        RECT 4.400 3.575 74.765 4.440 ;
  END
END CLA_16
END LIBRARY

