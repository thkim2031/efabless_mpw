magic
tech sky130B
magscale 1 2
timestamp 1661734572
<< obsli1 >>
rect 1104 2159 358892 397681
<< obsm1 >>
rect 750 8 358892 397712
<< metal2 >>
rect 3238 399200 3294 400000
rect 6366 399200 6422 400000
rect 9494 399200 9550 400000
rect 12622 399200 12678 400000
rect 15750 399200 15806 400000
rect 18878 399200 18934 400000
rect 22006 399200 22062 400000
rect 25134 399200 25190 400000
rect 28262 399200 28318 400000
rect 31390 399200 31446 400000
rect 34518 399200 34574 400000
rect 37646 399200 37702 400000
rect 40774 399200 40830 400000
rect 43902 399200 43958 400000
rect 47030 399200 47086 400000
rect 50158 399200 50214 400000
rect 53286 399200 53342 400000
rect 56414 399200 56470 400000
rect 59542 399200 59598 400000
rect 62670 399200 62726 400000
rect 65798 399200 65854 400000
rect 68926 399200 68982 400000
rect 72054 399200 72110 400000
rect 75182 399200 75238 400000
rect 78310 399200 78366 400000
rect 81438 399200 81494 400000
rect 84566 399200 84622 400000
rect 87694 399200 87750 400000
rect 90822 399200 90878 400000
rect 93950 399200 94006 400000
rect 97078 399200 97134 400000
rect 100206 399200 100262 400000
rect 103334 399200 103390 400000
rect 106462 399200 106518 400000
rect 109590 399200 109646 400000
rect 112718 399200 112774 400000
rect 115846 399200 115902 400000
rect 118974 399200 119030 400000
rect 122102 399200 122158 400000
rect 125230 399200 125286 400000
rect 128358 399200 128414 400000
rect 131486 399200 131542 400000
rect 134614 399200 134670 400000
rect 137742 399200 137798 400000
rect 140870 399200 140926 400000
rect 143998 399200 144054 400000
rect 147126 399200 147182 400000
rect 150254 399200 150310 400000
rect 153382 399200 153438 400000
rect 156510 399200 156566 400000
rect 159638 399200 159694 400000
rect 162766 399200 162822 400000
rect 165894 399200 165950 400000
rect 169022 399200 169078 400000
rect 172150 399200 172206 400000
rect 175278 399200 175334 400000
rect 178406 399200 178462 400000
rect 181534 399200 181590 400000
rect 184662 399200 184718 400000
rect 187790 399200 187846 400000
rect 190918 399200 190974 400000
rect 194046 399200 194102 400000
rect 197174 399200 197230 400000
rect 200302 399200 200358 400000
rect 203430 399200 203486 400000
rect 206558 399200 206614 400000
rect 209686 399200 209742 400000
rect 212814 399200 212870 400000
rect 215942 399200 215998 400000
rect 219070 399200 219126 400000
rect 222198 399200 222254 400000
rect 225326 399200 225382 400000
rect 228454 399200 228510 400000
rect 231582 399200 231638 400000
rect 234710 399200 234766 400000
rect 237838 399200 237894 400000
rect 240966 399200 241022 400000
rect 244094 399200 244150 400000
rect 247222 399200 247278 400000
rect 250350 399200 250406 400000
rect 253478 399200 253534 400000
rect 256606 399200 256662 400000
rect 259734 399200 259790 400000
rect 262862 399200 262918 400000
rect 265990 399200 266046 400000
rect 269118 399200 269174 400000
rect 272246 399200 272302 400000
rect 275374 399200 275430 400000
rect 278502 399200 278558 400000
rect 281630 399200 281686 400000
rect 284758 399200 284814 400000
rect 287886 399200 287942 400000
rect 291014 399200 291070 400000
rect 294142 399200 294198 400000
rect 297270 399200 297326 400000
rect 300398 399200 300454 400000
rect 303526 399200 303582 400000
rect 306654 399200 306710 400000
rect 309782 399200 309838 400000
rect 312910 399200 312966 400000
rect 316038 399200 316094 400000
rect 319166 399200 319222 400000
rect 322294 399200 322350 400000
rect 325422 399200 325478 400000
rect 328550 399200 328606 400000
rect 331678 399200 331734 400000
rect 334806 399200 334862 400000
rect 337934 399200 337990 400000
rect 341062 399200 341118 400000
rect 344190 399200 344246 400000
rect 347318 399200 347374 400000
rect 350446 399200 350502 400000
rect 353574 399200 353630 400000
rect 356702 399200 356758 400000
rect 21546 0 21602 800
rect 22190 0 22246 800
rect 22834 0 22890 800
rect 23478 0 23534 800
rect 24122 0 24178 800
rect 24766 0 24822 800
rect 25410 0 25466 800
rect 26054 0 26110 800
rect 26698 0 26754 800
rect 27342 0 27398 800
rect 27986 0 28042 800
rect 28630 0 28686 800
rect 29274 0 29330 800
rect 29918 0 29974 800
rect 30562 0 30618 800
rect 31206 0 31262 800
rect 31850 0 31906 800
rect 32494 0 32550 800
rect 33138 0 33194 800
rect 33782 0 33838 800
rect 34426 0 34482 800
rect 35070 0 35126 800
rect 35714 0 35770 800
rect 36358 0 36414 800
rect 37002 0 37058 800
rect 37646 0 37702 800
rect 38290 0 38346 800
rect 38934 0 38990 800
rect 39578 0 39634 800
rect 40222 0 40278 800
rect 40866 0 40922 800
rect 41510 0 41566 800
rect 42154 0 42210 800
rect 42798 0 42854 800
rect 43442 0 43498 800
rect 44086 0 44142 800
rect 44730 0 44786 800
rect 45374 0 45430 800
rect 46018 0 46074 800
rect 46662 0 46718 800
rect 47306 0 47362 800
rect 47950 0 48006 800
rect 48594 0 48650 800
rect 49238 0 49294 800
rect 49882 0 49938 800
rect 50526 0 50582 800
rect 51170 0 51226 800
rect 51814 0 51870 800
rect 52458 0 52514 800
rect 53102 0 53158 800
rect 53746 0 53802 800
rect 54390 0 54446 800
rect 55034 0 55090 800
rect 55678 0 55734 800
rect 56322 0 56378 800
rect 56966 0 57022 800
rect 57610 0 57666 800
rect 58254 0 58310 800
rect 58898 0 58954 800
rect 59542 0 59598 800
rect 60186 0 60242 800
rect 60830 0 60886 800
rect 61474 0 61530 800
rect 62118 0 62174 800
rect 62762 0 62818 800
rect 63406 0 63462 800
rect 64050 0 64106 800
rect 64694 0 64750 800
rect 65338 0 65394 800
rect 65982 0 66038 800
rect 66626 0 66682 800
rect 67270 0 67326 800
rect 67914 0 67970 800
rect 68558 0 68614 800
rect 69202 0 69258 800
rect 69846 0 69902 800
rect 70490 0 70546 800
rect 71134 0 71190 800
rect 71778 0 71834 800
rect 72422 0 72478 800
rect 73066 0 73122 800
rect 73710 0 73766 800
rect 74354 0 74410 800
rect 74998 0 75054 800
rect 75642 0 75698 800
rect 76286 0 76342 800
rect 76930 0 76986 800
rect 77574 0 77630 800
rect 78218 0 78274 800
rect 78862 0 78918 800
rect 79506 0 79562 800
rect 80150 0 80206 800
rect 80794 0 80850 800
rect 81438 0 81494 800
rect 82082 0 82138 800
rect 82726 0 82782 800
rect 83370 0 83426 800
rect 84014 0 84070 800
rect 84658 0 84714 800
rect 85302 0 85358 800
rect 85946 0 86002 800
rect 86590 0 86646 800
rect 87234 0 87290 800
rect 87878 0 87934 800
rect 88522 0 88578 800
rect 89166 0 89222 800
rect 89810 0 89866 800
rect 90454 0 90510 800
rect 91098 0 91154 800
rect 91742 0 91798 800
rect 92386 0 92442 800
rect 93030 0 93086 800
rect 93674 0 93730 800
rect 94318 0 94374 800
rect 94962 0 95018 800
rect 95606 0 95662 800
rect 96250 0 96306 800
rect 96894 0 96950 800
rect 97538 0 97594 800
rect 98182 0 98238 800
rect 98826 0 98882 800
rect 99470 0 99526 800
rect 100114 0 100170 800
rect 100758 0 100814 800
rect 101402 0 101458 800
rect 102046 0 102102 800
rect 102690 0 102746 800
rect 103334 0 103390 800
rect 103978 0 104034 800
rect 104622 0 104678 800
rect 105266 0 105322 800
rect 105910 0 105966 800
rect 106554 0 106610 800
rect 107198 0 107254 800
rect 107842 0 107898 800
rect 108486 0 108542 800
rect 109130 0 109186 800
rect 109774 0 109830 800
rect 110418 0 110474 800
rect 111062 0 111118 800
rect 111706 0 111762 800
rect 112350 0 112406 800
rect 112994 0 113050 800
rect 113638 0 113694 800
rect 114282 0 114338 800
rect 114926 0 114982 800
rect 115570 0 115626 800
rect 116214 0 116270 800
rect 116858 0 116914 800
rect 117502 0 117558 800
rect 118146 0 118202 800
rect 118790 0 118846 800
rect 119434 0 119490 800
rect 120078 0 120134 800
rect 120722 0 120778 800
rect 121366 0 121422 800
rect 122010 0 122066 800
rect 122654 0 122710 800
rect 123298 0 123354 800
rect 123942 0 123998 800
rect 124586 0 124642 800
rect 125230 0 125286 800
rect 125874 0 125930 800
rect 126518 0 126574 800
rect 127162 0 127218 800
rect 127806 0 127862 800
rect 128450 0 128506 800
rect 129094 0 129150 800
rect 129738 0 129794 800
rect 130382 0 130438 800
rect 131026 0 131082 800
rect 131670 0 131726 800
rect 132314 0 132370 800
rect 132958 0 133014 800
rect 133602 0 133658 800
rect 134246 0 134302 800
rect 134890 0 134946 800
rect 135534 0 135590 800
rect 136178 0 136234 800
rect 136822 0 136878 800
rect 137466 0 137522 800
rect 138110 0 138166 800
rect 138754 0 138810 800
rect 139398 0 139454 800
rect 140042 0 140098 800
rect 140686 0 140742 800
rect 141330 0 141386 800
rect 141974 0 142030 800
rect 142618 0 142674 800
rect 143262 0 143318 800
rect 143906 0 143962 800
rect 144550 0 144606 800
rect 145194 0 145250 800
rect 145838 0 145894 800
rect 146482 0 146538 800
rect 147126 0 147182 800
rect 147770 0 147826 800
rect 148414 0 148470 800
rect 149058 0 149114 800
rect 149702 0 149758 800
rect 150346 0 150402 800
rect 150990 0 151046 800
rect 151634 0 151690 800
rect 152278 0 152334 800
rect 152922 0 152978 800
rect 153566 0 153622 800
rect 154210 0 154266 800
rect 154854 0 154910 800
rect 155498 0 155554 800
rect 156142 0 156198 800
rect 156786 0 156842 800
rect 157430 0 157486 800
rect 158074 0 158130 800
rect 158718 0 158774 800
rect 159362 0 159418 800
rect 160006 0 160062 800
rect 160650 0 160706 800
rect 161294 0 161350 800
rect 161938 0 161994 800
rect 162582 0 162638 800
rect 163226 0 163282 800
rect 163870 0 163926 800
rect 164514 0 164570 800
rect 165158 0 165214 800
rect 165802 0 165858 800
rect 166446 0 166502 800
rect 167090 0 167146 800
rect 167734 0 167790 800
rect 168378 0 168434 800
rect 169022 0 169078 800
rect 169666 0 169722 800
rect 170310 0 170366 800
rect 170954 0 171010 800
rect 171598 0 171654 800
rect 172242 0 172298 800
rect 172886 0 172942 800
rect 173530 0 173586 800
rect 174174 0 174230 800
rect 174818 0 174874 800
rect 175462 0 175518 800
rect 176106 0 176162 800
rect 176750 0 176806 800
rect 177394 0 177450 800
rect 178038 0 178094 800
rect 178682 0 178738 800
rect 179326 0 179382 800
rect 179970 0 180026 800
rect 180614 0 180670 800
rect 181258 0 181314 800
rect 181902 0 181958 800
rect 182546 0 182602 800
rect 183190 0 183246 800
rect 183834 0 183890 800
rect 184478 0 184534 800
rect 185122 0 185178 800
rect 185766 0 185822 800
rect 186410 0 186466 800
rect 187054 0 187110 800
rect 187698 0 187754 800
rect 188342 0 188398 800
rect 188986 0 189042 800
rect 189630 0 189686 800
rect 190274 0 190330 800
rect 190918 0 190974 800
rect 191562 0 191618 800
rect 192206 0 192262 800
rect 192850 0 192906 800
rect 193494 0 193550 800
rect 194138 0 194194 800
rect 194782 0 194838 800
rect 195426 0 195482 800
rect 196070 0 196126 800
rect 196714 0 196770 800
rect 197358 0 197414 800
rect 198002 0 198058 800
rect 198646 0 198702 800
rect 199290 0 199346 800
rect 199934 0 199990 800
rect 200578 0 200634 800
rect 201222 0 201278 800
rect 201866 0 201922 800
rect 202510 0 202566 800
rect 203154 0 203210 800
rect 203798 0 203854 800
rect 204442 0 204498 800
rect 205086 0 205142 800
rect 205730 0 205786 800
rect 206374 0 206430 800
rect 207018 0 207074 800
rect 207662 0 207718 800
rect 208306 0 208362 800
rect 208950 0 209006 800
rect 209594 0 209650 800
rect 210238 0 210294 800
rect 210882 0 210938 800
rect 211526 0 211582 800
rect 212170 0 212226 800
rect 212814 0 212870 800
rect 213458 0 213514 800
rect 214102 0 214158 800
rect 214746 0 214802 800
rect 215390 0 215446 800
rect 216034 0 216090 800
rect 216678 0 216734 800
rect 217322 0 217378 800
rect 217966 0 218022 800
rect 218610 0 218666 800
rect 219254 0 219310 800
rect 219898 0 219954 800
rect 220542 0 220598 800
rect 221186 0 221242 800
rect 221830 0 221886 800
rect 222474 0 222530 800
rect 223118 0 223174 800
rect 223762 0 223818 800
rect 224406 0 224462 800
rect 225050 0 225106 800
rect 225694 0 225750 800
rect 226338 0 226394 800
rect 226982 0 227038 800
rect 227626 0 227682 800
rect 228270 0 228326 800
rect 228914 0 228970 800
rect 229558 0 229614 800
rect 230202 0 230258 800
rect 230846 0 230902 800
rect 231490 0 231546 800
rect 232134 0 232190 800
rect 232778 0 232834 800
rect 233422 0 233478 800
rect 234066 0 234122 800
rect 234710 0 234766 800
rect 235354 0 235410 800
rect 235998 0 236054 800
rect 236642 0 236698 800
rect 237286 0 237342 800
rect 237930 0 237986 800
rect 238574 0 238630 800
rect 239218 0 239274 800
rect 239862 0 239918 800
rect 240506 0 240562 800
rect 241150 0 241206 800
rect 241794 0 241850 800
rect 242438 0 242494 800
rect 243082 0 243138 800
rect 243726 0 243782 800
rect 244370 0 244426 800
rect 245014 0 245070 800
rect 245658 0 245714 800
rect 246302 0 246358 800
rect 246946 0 247002 800
rect 247590 0 247646 800
rect 248234 0 248290 800
rect 248878 0 248934 800
rect 249522 0 249578 800
rect 250166 0 250222 800
rect 250810 0 250866 800
rect 251454 0 251510 800
rect 252098 0 252154 800
rect 252742 0 252798 800
rect 253386 0 253442 800
rect 254030 0 254086 800
rect 254674 0 254730 800
rect 255318 0 255374 800
rect 255962 0 256018 800
rect 256606 0 256662 800
rect 257250 0 257306 800
rect 257894 0 257950 800
rect 258538 0 258594 800
rect 259182 0 259238 800
rect 259826 0 259882 800
rect 260470 0 260526 800
rect 261114 0 261170 800
rect 261758 0 261814 800
rect 262402 0 262458 800
rect 263046 0 263102 800
rect 263690 0 263746 800
rect 264334 0 264390 800
rect 264978 0 265034 800
rect 265622 0 265678 800
rect 266266 0 266322 800
rect 266910 0 266966 800
rect 267554 0 267610 800
rect 268198 0 268254 800
rect 268842 0 268898 800
rect 269486 0 269542 800
rect 270130 0 270186 800
rect 270774 0 270830 800
rect 271418 0 271474 800
rect 272062 0 272118 800
rect 272706 0 272762 800
rect 273350 0 273406 800
rect 273994 0 274050 800
rect 274638 0 274694 800
rect 275282 0 275338 800
rect 275926 0 275982 800
rect 276570 0 276626 800
rect 277214 0 277270 800
rect 277858 0 277914 800
rect 278502 0 278558 800
rect 279146 0 279202 800
rect 279790 0 279846 800
rect 280434 0 280490 800
rect 281078 0 281134 800
rect 281722 0 281778 800
rect 282366 0 282422 800
rect 283010 0 283066 800
rect 283654 0 283710 800
rect 284298 0 284354 800
rect 284942 0 284998 800
rect 285586 0 285642 800
rect 286230 0 286286 800
rect 286874 0 286930 800
rect 287518 0 287574 800
rect 288162 0 288218 800
rect 288806 0 288862 800
rect 289450 0 289506 800
rect 290094 0 290150 800
rect 290738 0 290794 800
rect 291382 0 291438 800
rect 292026 0 292082 800
rect 292670 0 292726 800
rect 293314 0 293370 800
rect 293958 0 294014 800
rect 294602 0 294658 800
rect 295246 0 295302 800
rect 295890 0 295946 800
rect 296534 0 296590 800
rect 297178 0 297234 800
rect 297822 0 297878 800
rect 298466 0 298522 800
rect 299110 0 299166 800
rect 299754 0 299810 800
rect 300398 0 300454 800
rect 301042 0 301098 800
rect 301686 0 301742 800
rect 302330 0 302386 800
rect 302974 0 303030 800
rect 303618 0 303674 800
rect 304262 0 304318 800
rect 304906 0 304962 800
rect 305550 0 305606 800
rect 306194 0 306250 800
rect 306838 0 306894 800
rect 307482 0 307538 800
rect 308126 0 308182 800
rect 308770 0 308826 800
rect 309414 0 309470 800
rect 310058 0 310114 800
rect 310702 0 310758 800
rect 311346 0 311402 800
rect 311990 0 312046 800
rect 312634 0 312690 800
rect 313278 0 313334 800
rect 313922 0 313978 800
rect 314566 0 314622 800
rect 315210 0 315266 800
rect 315854 0 315910 800
rect 316498 0 316554 800
rect 317142 0 317198 800
rect 317786 0 317842 800
rect 318430 0 318486 800
rect 319074 0 319130 800
rect 319718 0 319774 800
rect 320362 0 320418 800
rect 321006 0 321062 800
rect 321650 0 321706 800
rect 322294 0 322350 800
rect 322938 0 322994 800
rect 323582 0 323638 800
rect 324226 0 324282 800
rect 324870 0 324926 800
rect 325514 0 325570 800
rect 326158 0 326214 800
rect 326802 0 326858 800
rect 327446 0 327502 800
rect 328090 0 328146 800
rect 328734 0 328790 800
rect 329378 0 329434 800
rect 330022 0 330078 800
rect 330666 0 330722 800
rect 331310 0 331366 800
rect 331954 0 332010 800
rect 332598 0 332654 800
rect 333242 0 333298 800
rect 333886 0 333942 800
rect 334530 0 334586 800
rect 335174 0 335230 800
rect 335818 0 335874 800
rect 336462 0 336518 800
rect 337106 0 337162 800
rect 337750 0 337806 800
rect 338394 0 338450 800
<< obsm2 >>
rect 756 399144 3182 399200
rect 3350 399144 6310 399200
rect 6478 399144 9438 399200
rect 9606 399144 12566 399200
rect 12734 399144 15694 399200
rect 15862 399144 18822 399200
rect 18990 399144 21950 399200
rect 22118 399144 25078 399200
rect 25246 399144 28206 399200
rect 28374 399144 31334 399200
rect 31502 399144 34462 399200
rect 34630 399144 37590 399200
rect 37758 399144 40718 399200
rect 40886 399144 43846 399200
rect 44014 399144 46974 399200
rect 47142 399144 50102 399200
rect 50270 399144 53230 399200
rect 53398 399144 56358 399200
rect 56526 399144 59486 399200
rect 59654 399144 62614 399200
rect 62782 399144 65742 399200
rect 65910 399144 68870 399200
rect 69038 399144 71998 399200
rect 72166 399144 75126 399200
rect 75294 399144 78254 399200
rect 78422 399144 81382 399200
rect 81550 399144 84510 399200
rect 84678 399144 87638 399200
rect 87806 399144 90766 399200
rect 90934 399144 93894 399200
rect 94062 399144 97022 399200
rect 97190 399144 100150 399200
rect 100318 399144 103278 399200
rect 103446 399144 106406 399200
rect 106574 399144 109534 399200
rect 109702 399144 112662 399200
rect 112830 399144 115790 399200
rect 115958 399144 118918 399200
rect 119086 399144 122046 399200
rect 122214 399144 125174 399200
rect 125342 399144 128302 399200
rect 128470 399144 131430 399200
rect 131598 399144 134558 399200
rect 134726 399144 137686 399200
rect 137854 399144 140814 399200
rect 140982 399144 143942 399200
rect 144110 399144 147070 399200
rect 147238 399144 150198 399200
rect 150366 399144 153326 399200
rect 153494 399144 156454 399200
rect 156622 399144 159582 399200
rect 159750 399144 162710 399200
rect 162878 399144 165838 399200
rect 166006 399144 168966 399200
rect 169134 399144 172094 399200
rect 172262 399144 175222 399200
rect 175390 399144 178350 399200
rect 178518 399144 181478 399200
rect 181646 399144 184606 399200
rect 184774 399144 187734 399200
rect 187902 399144 190862 399200
rect 191030 399144 193990 399200
rect 194158 399144 197118 399200
rect 197286 399144 200246 399200
rect 200414 399144 203374 399200
rect 203542 399144 206502 399200
rect 206670 399144 209630 399200
rect 209798 399144 212758 399200
rect 212926 399144 215886 399200
rect 216054 399144 219014 399200
rect 219182 399144 222142 399200
rect 222310 399144 225270 399200
rect 225438 399144 228398 399200
rect 228566 399144 231526 399200
rect 231694 399144 234654 399200
rect 234822 399144 237782 399200
rect 237950 399144 240910 399200
rect 241078 399144 244038 399200
rect 244206 399144 247166 399200
rect 247334 399144 250294 399200
rect 250462 399144 253422 399200
rect 253590 399144 256550 399200
rect 256718 399144 259678 399200
rect 259846 399144 262806 399200
rect 262974 399144 265934 399200
rect 266102 399144 269062 399200
rect 269230 399144 272190 399200
rect 272358 399144 275318 399200
rect 275486 399144 278446 399200
rect 278614 399144 281574 399200
rect 281742 399144 284702 399200
rect 284870 399144 287830 399200
rect 287998 399144 290958 399200
rect 291126 399144 294086 399200
rect 294254 399144 297214 399200
rect 297382 399144 300342 399200
rect 300510 399144 303470 399200
rect 303638 399144 306598 399200
rect 306766 399144 309726 399200
rect 309894 399144 312854 399200
rect 313022 399144 315982 399200
rect 316150 399144 319110 399200
rect 319278 399144 322238 399200
rect 322406 399144 325366 399200
rect 325534 399144 328494 399200
rect 328662 399144 331622 399200
rect 331790 399144 334750 399200
rect 334918 399144 337878 399200
rect 338046 399144 341006 399200
rect 341174 399144 344134 399200
rect 344302 399144 347262 399200
rect 347430 399144 350390 399200
rect 350558 399144 353518 399200
rect 353686 399144 356646 399200
rect 356814 399144 357802 399200
rect 756 856 357802 399144
rect 756 2 21490 856
rect 21658 2 22134 856
rect 22302 2 22778 856
rect 22946 2 23422 856
rect 23590 2 24066 856
rect 24234 2 24710 856
rect 24878 2 25354 856
rect 25522 2 25998 856
rect 26166 2 26642 856
rect 26810 2 27286 856
rect 27454 2 27930 856
rect 28098 2 28574 856
rect 28742 2 29218 856
rect 29386 2 29862 856
rect 30030 2 30506 856
rect 30674 2 31150 856
rect 31318 2 31794 856
rect 31962 2 32438 856
rect 32606 2 33082 856
rect 33250 2 33726 856
rect 33894 2 34370 856
rect 34538 2 35014 856
rect 35182 2 35658 856
rect 35826 2 36302 856
rect 36470 2 36946 856
rect 37114 2 37590 856
rect 37758 2 38234 856
rect 38402 2 38878 856
rect 39046 2 39522 856
rect 39690 2 40166 856
rect 40334 2 40810 856
rect 40978 2 41454 856
rect 41622 2 42098 856
rect 42266 2 42742 856
rect 42910 2 43386 856
rect 43554 2 44030 856
rect 44198 2 44674 856
rect 44842 2 45318 856
rect 45486 2 45962 856
rect 46130 2 46606 856
rect 46774 2 47250 856
rect 47418 2 47894 856
rect 48062 2 48538 856
rect 48706 2 49182 856
rect 49350 2 49826 856
rect 49994 2 50470 856
rect 50638 2 51114 856
rect 51282 2 51758 856
rect 51926 2 52402 856
rect 52570 2 53046 856
rect 53214 2 53690 856
rect 53858 2 54334 856
rect 54502 2 54978 856
rect 55146 2 55622 856
rect 55790 2 56266 856
rect 56434 2 56910 856
rect 57078 2 57554 856
rect 57722 2 58198 856
rect 58366 2 58842 856
rect 59010 2 59486 856
rect 59654 2 60130 856
rect 60298 2 60774 856
rect 60942 2 61418 856
rect 61586 2 62062 856
rect 62230 2 62706 856
rect 62874 2 63350 856
rect 63518 2 63994 856
rect 64162 2 64638 856
rect 64806 2 65282 856
rect 65450 2 65926 856
rect 66094 2 66570 856
rect 66738 2 67214 856
rect 67382 2 67858 856
rect 68026 2 68502 856
rect 68670 2 69146 856
rect 69314 2 69790 856
rect 69958 2 70434 856
rect 70602 2 71078 856
rect 71246 2 71722 856
rect 71890 2 72366 856
rect 72534 2 73010 856
rect 73178 2 73654 856
rect 73822 2 74298 856
rect 74466 2 74942 856
rect 75110 2 75586 856
rect 75754 2 76230 856
rect 76398 2 76874 856
rect 77042 2 77518 856
rect 77686 2 78162 856
rect 78330 2 78806 856
rect 78974 2 79450 856
rect 79618 2 80094 856
rect 80262 2 80738 856
rect 80906 2 81382 856
rect 81550 2 82026 856
rect 82194 2 82670 856
rect 82838 2 83314 856
rect 83482 2 83958 856
rect 84126 2 84602 856
rect 84770 2 85246 856
rect 85414 2 85890 856
rect 86058 2 86534 856
rect 86702 2 87178 856
rect 87346 2 87822 856
rect 87990 2 88466 856
rect 88634 2 89110 856
rect 89278 2 89754 856
rect 89922 2 90398 856
rect 90566 2 91042 856
rect 91210 2 91686 856
rect 91854 2 92330 856
rect 92498 2 92974 856
rect 93142 2 93618 856
rect 93786 2 94262 856
rect 94430 2 94906 856
rect 95074 2 95550 856
rect 95718 2 96194 856
rect 96362 2 96838 856
rect 97006 2 97482 856
rect 97650 2 98126 856
rect 98294 2 98770 856
rect 98938 2 99414 856
rect 99582 2 100058 856
rect 100226 2 100702 856
rect 100870 2 101346 856
rect 101514 2 101990 856
rect 102158 2 102634 856
rect 102802 2 103278 856
rect 103446 2 103922 856
rect 104090 2 104566 856
rect 104734 2 105210 856
rect 105378 2 105854 856
rect 106022 2 106498 856
rect 106666 2 107142 856
rect 107310 2 107786 856
rect 107954 2 108430 856
rect 108598 2 109074 856
rect 109242 2 109718 856
rect 109886 2 110362 856
rect 110530 2 111006 856
rect 111174 2 111650 856
rect 111818 2 112294 856
rect 112462 2 112938 856
rect 113106 2 113582 856
rect 113750 2 114226 856
rect 114394 2 114870 856
rect 115038 2 115514 856
rect 115682 2 116158 856
rect 116326 2 116802 856
rect 116970 2 117446 856
rect 117614 2 118090 856
rect 118258 2 118734 856
rect 118902 2 119378 856
rect 119546 2 120022 856
rect 120190 2 120666 856
rect 120834 2 121310 856
rect 121478 2 121954 856
rect 122122 2 122598 856
rect 122766 2 123242 856
rect 123410 2 123886 856
rect 124054 2 124530 856
rect 124698 2 125174 856
rect 125342 2 125818 856
rect 125986 2 126462 856
rect 126630 2 127106 856
rect 127274 2 127750 856
rect 127918 2 128394 856
rect 128562 2 129038 856
rect 129206 2 129682 856
rect 129850 2 130326 856
rect 130494 2 130970 856
rect 131138 2 131614 856
rect 131782 2 132258 856
rect 132426 2 132902 856
rect 133070 2 133546 856
rect 133714 2 134190 856
rect 134358 2 134834 856
rect 135002 2 135478 856
rect 135646 2 136122 856
rect 136290 2 136766 856
rect 136934 2 137410 856
rect 137578 2 138054 856
rect 138222 2 138698 856
rect 138866 2 139342 856
rect 139510 2 139986 856
rect 140154 2 140630 856
rect 140798 2 141274 856
rect 141442 2 141918 856
rect 142086 2 142562 856
rect 142730 2 143206 856
rect 143374 2 143850 856
rect 144018 2 144494 856
rect 144662 2 145138 856
rect 145306 2 145782 856
rect 145950 2 146426 856
rect 146594 2 147070 856
rect 147238 2 147714 856
rect 147882 2 148358 856
rect 148526 2 149002 856
rect 149170 2 149646 856
rect 149814 2 150290 856
rect 150458 2 150934 856
rect 151102 2 151578 856
rect 151746 2 152222 856
rect 152390 2 152866 856
rect 153034 2 153510 856
rect 153678 2 154154 856
rect 154322 2 154798 856
rect 154966 2 155442 856
rect 155610 2 156086 856
rect 156254 2 156730 856
rect 156898 2 157374 856
rect 157542 2 158018 856
rect 158186 2 158662 856
rect 158830 2 159306 856
rect 159474 2 159950 856
rect 160118 2 160594 856
rect 160762 2 161238 856
rect 161406 2 161882 856
rect 162050 2 162526 856
rect 162694 2 163170 856
rect 163338 2 163814 856
rect 163982 2 164458 856
rect 164626 2 165102 856
rect 165270 2 165746 856
rect 165914 2 166390 856
rect 166558 2 167034 856
rect 167202 2 167678 856
rect 167846 2 168322 856
rect 168490 2 168966 856
rect 169134 2 169610 856
rect 169778 2 170254 856
rect 170422 2 170898 856
rect 171066 2 171542 856
rect 171710 2 172186 856
rect 172354 2 172830 856
rect 172998 2 173474 856
rect 173642 2 174118 856
rect 174286 2 174762 856
rect 174930 2 175406 856
rect 175574 2 176050 856
rect 176218 2 176694 856
rect 176862 2 177338 856
rect 177506 2 177982 856
rect 178150 2 178626 856
rect 178794 2 179270 856
rect 179438 2 179914 856
rect 180082 2 180558 856
rect 180726 2 181202 856
rect 181370 2 181846 856
rect 182014 2 182490 856
rect 182658 2 183134 856
rect 183302 2 183778 856
rect 183946 2 184422 856
rect 184590 2 185066 856
rect 185234 2 185710 856
rect 185878 2 186354 856
rect 186522 2 186998 856
rect 187166 2 187642 856
rect 187810 2 188286 856
rect 188454 2 188930 856
rect 189098 2 189574 856
rect 189742 2 190218 856
rect 190386 2 190862 856
rect 191030 2 191506 856
rect 191674 2 192150 856
rect 192318 2 192794 856
rect 192962 2 193438 856
rect 193606 2 194082 856
rect 194250 2 194726 856
rect 194894 2 195370 856
rect 195538 2 196014 856
rect 196182 2 196658 856
rect 196826 2 197302 856
rect 197470 2 197946 856
rect 198114 2 198590 856
rect 198758 2 199234 856
rect 199402 2 199878 856
rect 200046 2 200522 856
rect 200690 2 201166 856
rect 201334 2 201810 856
rect 201978 2 202454 856
rect 202622 2 203098 856
rect 203266 2 203742 856
rect 203910 2 204386 856
rect 204554 2 205030 856
rect 205198 2 205674 856
rect 205842 2 206318 856
rect 206486 2 206962 856
rect 207130 2 207606 856
rect 207774 2 208250 856
rect 208418 2 208894 856
rect 209062 2 209538 856
rect 209706 2 210182 856
rect 210350 2 210826 856
rect 210994 2 211470 856
rect 211638 2 212114 856
rect 212282 2 212758 856
rect 212926 2 213402 856
rect 213570 2 214046 856
rect 214214 2 214690 856
rect 214858 2 215334 856
rect 215502 2 215978 856
rect 216146 2 216622 856
rect 216790 2 217266 856
rect 217434 2 217910 856
rect 218078 2 218554 856
rect 218722 2 219198 856
rect 219366 2 219842 856
rect 220010 2 220486 856
rect 220654 2 221130 856
rect 221298 2 221774 856
rect 221942 2 222418 856
rect 222586 2 223062 856
rect 223230 2 223706 856
rect 223874 2 224350 856
rect 224518 2 224994 856
rect 225162 2 225638 856
rect 225806 2 226282 856
rect 226450 2 226926 856
rect 227094 2 227570 856
rect 227738 2 228214 856
rect 228382 2 228858 856
rect 229026 2 229502 856
rect 229670 2 230146 856
rect 230314 2 230790 856
rect 230958 2 231434 856
rect 231602 2 232078 856
rect 232246 2 232722 856
rect 232890 2 233366 856
rect 233534 2 234010 856
rect 234178 2 234654 856
rect 234822 2 235298 856
rect 235466 2 235942 856
rect 236110 2 236586 856
rect 236754 2 237230 856
rect 237398 2 237874 856
rect 238042 2 238518 856
rect 238686 2 239162 856
rect 239330 2 239806 856
rect 239974 2 240450 856
rect 240618 2 241094 856
rect 241262 2 241738 856
rect 241906 2 242382 856
rect 242550 2 243026 856
rect 243194 2 243670 856
rect 243838 2 244314 856
rect 244482 2 244958 856
rect 245126 2 245602 856
rect 245770 2 246246 856
rect 246414 2 246890 856
rect 247058 2 247534 856
rect 247702 2 248178 856
rect 248346 2 248822 856
rect 248990 2 249466 856
rect 249634 2 250110 856
rect 250278 2 250754 856
rect 250922 2 251398 856
rect 251566 2 252042 856
rect 252210 2 252686 856
rect 252854 2 253330 856
rect 253498 2 253974 856
rect 254142 2 254618 856
rect 254786 2 255262 856
rect 255430 2 255906 856
rect 256074 2 256550 856
rect 256718 2 257194 856
rect 257362 2 257838 856
rect 258006 2 258482 856
rect 258650 2 259126 856
rect 259294 2 259770 856
rect 259938 2 260414 856
rect 260582 2 261058 856
rect 261226 2 261702 856
rect 261870 2 262346 856
rect 262514 2 262990 856
rect 263158 2 263634 856
rect 263802 2 264278 856
rect 264446 2 264922 856
rect 265090 2 265566 856
rect 265734 2 266210 856
rect 266378 2 266854 856
rect 267022 2 267498 856
rect 267666 2 268142 856
rect 268310 2 268786 856
rect 268954 2 269430 856
rect 269598 2 270074 856
rect 270242 2 270718 856
rect 270886 2 271362 856
rect 271530 2 272006 856
rect 272174 2 272650 856
rect 272818 2 273294 856
rect 273462 2 273938 856
rect 274106 2 274582 856
rect 274750 2 275226 856
rect 275394 2 275870 856
rect 276038 2 276514 856
rect 276682 2 277158 856
rect 277326 2 277802 856
rect 277970 2 278446 856
rect 278614 2 279090 856
rect 279258 2 279734 856
rect 279902 2 280378 856
rect 280546 2 281022 856
rect 281190 2 281666 856
rect 281834 2 282310 856
rect 282478 2 282954 856
rect 283122 2 283598 856
rect 283766 2 284242 856
rect 284410 2 284886 856
rect 285054 2 285530 856
rect 285698 2 286174 856
rect 286342 2 286818 856
rect 286986 2 287462 856
rect 287630 2 288106 856
rect 288274 2 288750 856
rect 288918 2 289394 856
rect 289562 2 290038 856
rect 290206 2 290682 856
rect 290850 2 291326 856
rect 291494 2 291970 856
rect 292138 2 292614 856
rect 292782 2 293258 856
rect 293426 2 293902 856
rect 294070 2 294546 856
rect 294714 2 295190 856
rect 295358 2 295834 856
rect 296002 2 296478 856
rect 296646 2 297122 856
rect 297290 2 297766 856
rect 297934 2 298410 856
rect 298578 2 299054 856
rect 299222 2 299698 856
rect 299866 2 300342 856
rect 300510 2 300986 856
rect 301154 2 301630 856
rect 301798 2 302274 856
rect 302442 2 302918 856
rect 303086 2 303562 856
rect 303730 2 304206 856
rect 304374 2 304850 856
rect 305018 2 305494 856
rect 305662 2 306138 856
rect 306306 2 306782 856
rect 306950 2 307426 856
rect 307594 2 308070 856
rect 308238 2 308714 856
rect 308882 2 309358 856
rect 309526 2 310002 856
rect 310170 2 310646 856
rect 310814 2 311290 856
rect 311458 2 311934 856
rect 312102 2 312578 856
rect 312746 2 313222 856
rect 313390 2 313866 856
rect 314034 2 314510 856
rect 314678 2 315154 856
rect 315322 2 315798 856
rect 315966 2 316442 856
rect 316610 2 317086 856
rect 317254 2 317730 856
rect 317898 2 318374 856
rect 318542 2 319018 856
rect 319186 2 319662 856
rect 319830 2 320306 856
rect 320474 2 320950 856
rect 321118 2 321594 856
rect 321762 2 322238 856
rect 322406 2 322882 856
rect 323050 2 323526 856
rect 323694 2 324170 856
rect 324338 2 324814 856
rect 324982 2 325458 856
rect 325626 2 326102 856
rect 326270 2 326746 856
rect 326914 2 327390 856
rect 327558 2 328034 856
rect 328202 2 328678 856
rect 328846 2 329322 856
rect 329490 2 329966 856
rect 330134 2 330610 856
rect 330778 2 331254 856
rect 331422 2 331898 856
rect 332066 2 332542 856
rect 332710 2 333186 856
rect 333354 2 333830 856
rect 333998 2 334474 856
rect 334642 2 335118 856
rect 335286 2 335762 856
rect 335930 2 336406 856
rect 336574 2 337050 856
rect 337218 2 337694 856
rect 337862 2 338338 856
rect 338506 2 357802 856
<< obsm3 >>
rect 1025 1123 357806 397697
<< metal4 >>
rect -1076 -4 -756 399844
rect -416 656 -96 399184
rect 4208 260614 4528 399844
rect 19568 260614 19888 399844
rect 34928 260614 35248 399844
rect 50288 260614 50608 399844
rect 65648 260614 65968 399844
rect 81008 260614 81328 399844
rect 96368 260614 96688 399844
rect 111728 260614 112048 399844
rect 4208 122410 4528 138000
rect 19568 122410 19888 138000
rect 34928 122410 35248 138000
rect 50288 122410 50608 138000
rect 65648 122410 65968 138000
rect 81008 122410 81328 138000
rect 96368 122410 96688 138000
rect 111728 122410 112048 138000
rect 127088 -4 127408 399844
rect 142448 304463 142768 399844
rect 157808 304463 158128 399844
rect 173168 304463 173488 399844
rect 188528 304463 188848 399844
rect 203888 304463 204208 399844
rect 219248 304463 219568 399844
rect 234608 304463 234928 399844
rect 249968 304463 250288 399844
rect 265328 304463 265648 399844
rect 280688 304463 281008 399844
rect 296048 304463 296368 399844
rect 129100 137040 129420 261168
rect 127996 2128 128316 88176
rect 142448 87428 142768 138000
rect 157808 87428 158128 138000
rect 173168 87428 173488 138000
rect 188528 87428 188848 138000
rect 203888 87428 204208 138000
rect 219248 87428 219568 138000
rect 234608 -4 234928 138000
rect 249968 -4 250288 138000
rect 265328 -4 265648 138000
rect 280688 -4 281008 138000
rect 296048 -4 296368 138000
rect 311408 -4 311728 399844
rect 326768 -4 327088 399844
rect 342128 -4 342448 399844
rect 357488 -4 357808 399844
rect 360092 656 360412 399184
rect 360752 -4 361072 399844
<< obsm4 >>
rect 1347 260534 4128 299984
rect 4608 260534 19488 299984
rect 19968 260534 34848 299984
rect 35328 260534 50208 299984
rect 50688 260534 65568 299984
rect 66048 260534 80928 299984
rect 81408 260534 96288 299984
rect 96768 260534 111648 299984
rect 112128 260534 127008 299984
rect 1347 138080 127008 260534
rect 1347 122330 4128 138080
rect 4608 122330 19488 138080
rect 19968 122330 34848 138080
rect 35328 122330 50208 138080
rect 50688 122330 65568 138080
rect 66048 122330 80928 138080
rect 81408 122330 96288 138080
rect 96768 122330 111648 138080
rect 112128 122330 127008 138080
rect 1347 1259 127008 122330
rect 127488 261248 298128 299984
rect 127488 136960 129020 261248
rect 129500 138080 298128 261248
rect 129500 136960 142368 138080
rect 127488 88256 142368 136960
rect 127488 2048 127916 88256
rect 128396 87348 142368 88256
rect 142848 87348 157728 138080
rect 158208 87348 173088 138080
rect 173568 87348 188448 138080
rect 188928 87348 203808 138080
rect 204288 87348 219168 138080
rect 219648 87348 234528 138080
rect 128396 2048 234528 87348
rect 127488 1259 234528 2048
rect 235008 1259 249888 138080
rect 250368 1259 265248 138080
rect 265728 1259 280608 138080
rect 281088 1259 295968 138080
rect 296448 1259 298128 138080
<< metal5 >>
rect -1076 399524 361072 399844
rect -416 398864 360412 399184
rect -1076 388296 361072 388616
rect -1076 372978 361072 373298
rect -1076 357660 361072 357980
rect -1076 342342 361072 342662
rect -1076 327024 361072 327344
rect -1076 311706 361072 312026
rect -1076 296388 361072 296708
rect -1076 281070 361072 281390
rect -1076 265752 361072 266072
rect -1076 250434 361072 250754
rect -1076 235116 361072 235436
rect -1076 219798 361072 220118
rect -1076 204480 361072 204800
rect -1076 189162 361072 189482
rect -1076 173844 361072 174164
rect -1076 158526 361072 158846
rect -1076 143208 361072 143528
rect 1056 130060 142768 130380
rect -1076 127890 361072 128210
rect -1076 112572 361072 112892
rect -1076 97254 361072 97574
rect -1076 81936 361072 82256
rect -1076 66618 361072 66938
rect -1076 51300 361072 51620
rect -1076 35982 361072 36302
rect -1076 20664 361072 20984
rect -1076 5346 361072 5666
rect -416 656 360412 976
rect -1076 -4 361072 316
<< labels >>
rlabel metal2 s 3238 399200 3294 400000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 97078 399200 97134 400000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 106462 399200 106518 400000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 115846 399200 115902 400000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 125230 399200 125286 400000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 134614 399200 134670 400000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 143998 399200 144054 400000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 153382 399200 153438 400000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 162766 399200 162822 400000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 172150 399200 172206 400000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 181534 399200 181590 400000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 12622 399200 12678 400000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 190918 399200 190974 400000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 200302 399200 200358 400000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 209686 399200 209742 400000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 219070 399200 219126 400000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 228454 399200 228510 400000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 237838 399200 237894 400000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 247222 399200 247278 400000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 256606 399200 256662 400000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 265990 399200 266046 400000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 275374 399200 275430 400000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 22006 399200 22062 400000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 284758 399200 284814 400000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 294142 399200 294198 400000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 303526 399200 303582 400000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 312910 399200 312966 400000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 322294 399200 322350 400000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 331678 399200 331734 400000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 341062 399200 341118 400000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 350446 399200 350502 400000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 31390 399200 31446 400000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 40774 399200 40830 400000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 50158 399200 50214 400000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 59542 399200 59598 400000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 68926 399200 68982 400000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 78310 399200 78366 400000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 87694 399200 87750 400000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6366 399200 6422 400000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 100206 399200 100262 400000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 109590 399200 109646 400000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 118974 399200 119030 400000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 128358 399200 128414 400000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 137742 399200 137798 400000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 147126 399200 147182 400000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 156510 399200 156566 400000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 165894 399200 165950 400000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 175278 399200 175334 400000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 184662 399200 184718 400000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 15750 399200 15806 400000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 194046 399200 194102 400000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 203430 399200 203486 400000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 212814 399200 212870 400000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 222198 399200 222254 400000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 231582 399200 231638 400000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 240966 399200 241022 400000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 250350 399200 250406 400000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 259734 399200 259790 400000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 269118 399200 269174 400000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 278502 399200 278558 400000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 25134 399200 25190 400000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 287886 399200 287942 400000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 297270 399200 297326 400000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 306654 399200 306710 400000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 316038 399200 316094 400000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 325422 399200 325478 400000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 334806 399200 334862 400000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 344190 399200 344246 400000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 353574 399200 353630 400000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 34518 399200 34574 400000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 43902 399200 43958 400000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 53286 399200 53342 400000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 62670 399200 62726 400000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 72054 399200 72110 400000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 81438 399200 81494 400000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 90822 399200 90878 400000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 9494 399200 9550 400000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 103334 399200 103390 400000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 112718 399200 112774 400000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 122102 399200 122158 400000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 131486 399200 131542 400000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 140870 399200 140926 400000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 150254 399200 150310 400000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 159638 399200 159694 400000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 169022 399200 169078 400000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 178406 399200 178462 400000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 187790 399200 187846 400000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 18878 399200 18934 400000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 197174 399200 197230 400000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 206558 399200 206614 400000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 215942 399200 215998 400000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 225326 399200 225382 400000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 234710 399200 234766 400000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 244094 399200 244150 400000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 253478 399200 253534 400000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 262862 399200 262918 400000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 272246 399200 272302 400000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 281630 399200 281686 400000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 28262 399200 28318 400000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 291014 399200 291070 400000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 300398 399200 300454 400000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 309782 399200 309838 400000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 319166 399200 319222 400000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 328550 399200 328606 400000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 337934 399200 337990 400000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 347318 399200 347374 400000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 356702 399200 356758 400000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 37646 399200 37702 400000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 47030 399200 47086 400000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 56414 399200 56470 400000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 65798 399200 65854 400000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 75182 399200 75238 400000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 84566 399200 84622 400000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 93950 399200 94006 400000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 337106 0 337162 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 337750 0 337806 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 338394 0 338450 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 89810 0 89866 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 283010 0 283066 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 284942 0 284998 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 286874 0 286930 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 288806 0 288862 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 290738 0 290794 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 292670 0 292726 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 294602 0 294658 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 296534 0 296590 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 298466 0 298522 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 300398 0 300454 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 302330 0 302386 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 304262 0 304318 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 306194 0 306250 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 308126 0 308182 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 310058 0 310114 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 311990 0 312046 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 313922 0 313978 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 315854 0 315910 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 317786 0 317842 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 319718 0 319774 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 111062 0 111118 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 321650 0 321706 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 323582 0 323638 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 325514 0 325570 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 327446 0 327502 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 329378 0 329434 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 331310 0 331366 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 333242 0 333298 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 335174 0 335230 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 114926 0 114982 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 118790 0 118846 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 120722 0 120778 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 124586 0 124642 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 128450 0 128506 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 132314 0 132370 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 93674 0 93730 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 147770 0 147826 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 149702 0 149758 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 153566 0 153622 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 159362 0 159418 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 163226 0 163282 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 167090 0 167146 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 170954 0 171010 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 178682 0 178738 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 180614 0 180670 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 182546 0 182602 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 184478 0 184534 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 97538 0 97594 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 186410 0 186466 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 188342 0 188398 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 190274 0 190330 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 192206 0 192262 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 196070 0 196126 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 198002 0 198058 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 199934 0 199990 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 201866 0 201922 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 203798 0 203854 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 99470 0 99526 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 205730 0 205786 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 207662 0 207718 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 209594 0 209650 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 211526 0 211582 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 213458 0 213514 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 217322 0 217378 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 219254 0 219310 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 221186 0 221242 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 223118 0 223174 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 101402 0 101458 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 225050 0 225106 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 226982 0 227038 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 228914 0 228970 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 230846 0 230902 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 232778 0 232834 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 234710 0 234766 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 238574 0 238630 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 240506 0 240562 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 242438 0 242494 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 103334 0 103390 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 244370 0 244426 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 246302 0 246358 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 250166 0 250222 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 252098 0 252154 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 254030 0 254086 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 255962 0 256018 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 257894 0 257950 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 259826 0 259882 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 261758 0 261814 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 105266 0 105322 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 263690 0 263746 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 265622 0 265678 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 267554 0 267610 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 269486 0 269542 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 271418 0 271474 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 273350 0 273406 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 275282 0 275338 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 277214 0 277270 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 279146 0 279202 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 281078 0 281134 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 107198 0 107254 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 283654 0 283710 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 285586 0 285642 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 287518 0 287574 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 289450 0 289506 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 291382 0 291438 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 293314 0 293370 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 295246 0 295302 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 297178 0 297234 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 299110 0 299166 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 301042 0 301098 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 109774 0 109830 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 302974 0 303030 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 304906 0 304962 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 306838 0 306894 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 308770 0 308826 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 310702 0 310758 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 312634 0 312690 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 314566 0 314622 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 316498 0 316554 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 318430 0 318486 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 320362 0 320418 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 111706 0 111762 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 322294 0 322350 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 324226 0 324282 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 326158 0 326214 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 328090 0 328146 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 330022 0 330078 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 331954 0 332010 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 333886 0 333942 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 335818 0 335874 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 113638 0 113694 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 121366 0 121422 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 123298 0 123354 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 125230 0 125286 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 127162 0 127218 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 92386 0 92442 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 129094 0 129150 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 132958 0 133014 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 134890 0 134946 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 136822 0 136878 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 138754 0 138810 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 140686 0 140742 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 142618 0 142674 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 144550 0 144606 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 150346 0 150402 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 154210 0 154266 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 158074 0 158130 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 160006 0 160062 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 161938 0 161994 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 96250 0 96306 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 167734 0 167790 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 169666 0 169722 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 171598 0 171654 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 173530 0 173586 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 175462 0 175518 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 177394 0 177450 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 181258 0 181314 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 185122 0 185178 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 98182 0 98238 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 187054 0 187110 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 188986 0 189042 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 190918 0 190974 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 192850 0 192906 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 194782 0 194838 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 196714 0 196770 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 198646 0 198702 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 200578 0 200634 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 202510 0 202566 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 204442 0 204498 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 206374 0 206430 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 208306 0 208362 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 210238 0 210294 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 212170 0 212226 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 214102 0 214158 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 216034 0 216090 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 217966 0 218022 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 219898 0 219954 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 221830 0 221886 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 223762 0 223818 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 225694 0 225750 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 227626 0 227682 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 229558 0 229614 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 231490 0 231546 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 233422 0 233478 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 235354 0 235410 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 237286 0 237342 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 239218 0 239274 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 241150 0 241206 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 243082 0 243138 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 245014 0 245070 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 246946 0 247002 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 248878 0 248934 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 250810 0 250866 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 252742 0 252798 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 254674 0 254730 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 256606 0 256662 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 258538 0 258594 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 262402 0 262458 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 105910 0 105966 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 264334 0 264390 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 266266 0 266322 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 268198 0 268254 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 270130 0 270186 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 272062 0 272118 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 273994 0 274050 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 275926 0 275982 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 279790 0 279846 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 281722 0 281778 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 91098 0 91154 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 284298 0 284354 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 286230 0 286286 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 288162 0 288218 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 290094 0 290150 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 292026 0 292082 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 293958 0 294014 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 295890 0 295946 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 297822 0 297878 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 299754 0 299810 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 301686 0 301742 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 110418 0 110474 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 303618 0 303674 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 305550 0 305606 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 307482 0 307538 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 309414 0 309470 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 311346 0 311402 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 313278 0 313334 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 315210 0 315266 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 317142 0 317198 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 319074 0 319130 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 321006 0 321062 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 322938 0 322994 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 324870 0 324926 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 326802 0 326858 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 328734 0 328790 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 330666 0 330722 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 332598 0 332654 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 334530 0 334586 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 336462 0 336518 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 116214 0 116270 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 120078 0 120134 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 123942 0 123998 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 127806 0 127862 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 133602 0 133658 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 141330 0 141386 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 94962 0 95018 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 156786 0 156842 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 164514 0 164570 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 96894 0 96950 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 168378 0 168434 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 172242 0 172298 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 176106 0 176162 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 179970 0 180026 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 181902 0 181958 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 183834 0 183890 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 185766 0 185822 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 98826 0 98882 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 187698 0 187754 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 189630 0 189686 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 191562 0 191618 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 193494 0 193550 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 195426 0 195482 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 197358 0 197414 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 199290 0 199346 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 201222 0 201278 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 203154 0 203210 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 205086 0 205142 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 207018 0 207074 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 208950 0 209006 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 210882 0 210938 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 212814 0 212870 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 214746 0 214802 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 216678 0 216734 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 218610 0 218666 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 220542 0 220598 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 222474 0 222530 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 224406 0 224462 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 102690 0 102746 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 226338 0 226394 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 228270 0 228326 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 230202 0 230258 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 232134 0 232190 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 234066 0 234122 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 235998 0 236054 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 237930 0 237986 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 239862 0 239918 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 241794 0 241850 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 243726 0 243782 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 245658 0 245714 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 247590 0 247646 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 249522 0 249578 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 251454 0 251510 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 253386 0 253442 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 255318 0 255374 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 257250 0 257306 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 259182 0 259238 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 261114 0 261170 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 263046 0 263102 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 106554 0 106610 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 264978 0 265034 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 266910 0 266966 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 268842 0 268898 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 270774 0 270830 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 272706 0 272762 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 274638 0 274694 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 276570 0 276626 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 278502 0 278558 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 280434 0 280490 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 282366 0 282422 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s -416 656 -96 399184 4 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -416 656 360412 976 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -416 398864 360412 399184 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 360092 656 360412 399184 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 4208 122410 4528 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 4208 260614 4528 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 122410 35248 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 34928 260614 35248 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 122410 65968 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 65648 260614 65968 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 122410 96688 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 96368 260614 96688 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 127088 -4 127408 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 87428 158128 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 157808 304463 158128 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 87428 188848 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 188528 304463 188848 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 87428 219568 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 219248 304463 219568 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 -4 250288 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 249968 304463 250288 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 -4 281008 138000 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 280688 304463 281008 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 311408 -4 311728 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s 342128 -4 342448 399844 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 5346 361072 5666 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 35982 361072 36302 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 66618 361072 66938 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 97254 361072 97574 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 127890 361072 128210 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 158526 361072 158846 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 189162 361072 189482 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 219798 361072 220118 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 250434 361072 250754 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 281070 361072 281390 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 311706 361072 312026 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 342342 361072 342662 6 vccd1
port 502 nsew power bidirectional
rlabel metal5 s -1076 372978 361072 373298 6 vccd1
port 502 nsew power bidirectional
rlabel metal4 s -1076 -4 -756 399844 4 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 -4 361072 316 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 399524 361072 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 360752 -4 361072 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 19568 122410 19888 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 19568 260614 19888 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 122410 50608 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 50288 260614 50608 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 122410 81328 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 81008 260614 81328 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 122410 112048 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 111728 260614 112048 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 87428 142768 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 142448 304463 142768 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 87428 173488 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 173168 304463 173488 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 87428 204208 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 203888 304463 204208 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 -4 234928 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 234608 304463 234928 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 -4 265648 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 265328 304463 265648 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 -4 296368 138000 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 296048 304463 296368 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 326768 -4 327088 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 357488 -4 357808 399844 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 20664 361072 20984 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 51300 361072 51620 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 81936 361072 82256 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 112572 361072 112892 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 143208 361072 143528 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 173844 361072 174164 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 204480 361072 204800 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 235116 361072 235436 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 265752 361072 266072 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 296388 361072 296708 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 327024 361072 327344 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 357660 361072 357980 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s -1076 388296 361072 388616 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 127996 2128 128316 88176 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 129100 137040 129420 261168 6 vssd1
port 503 nsew ground bidirectional
rlabel metal5 s 1056 130060 142768 130380 6 vssd1
port 503 nsew ground bidirectional
rlabel metal2 s 21546 0 21602 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 25410 0 25466 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 51170 0 51226 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 60830 0 60886 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 68558 0 68614 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 72422 0 72478 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 74354 0 74410 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 76286 0 76342 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 80150 0 80206 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 85946 0 86002 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 35714 0 35770 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 43442 0 43498 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 23478 0 23534 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 49882 0 49938 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 55678 0 55734 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 67270 0 67326 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 69202 0 69258 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 71134 0 71190 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 76930 0 76986 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 78862 0 78918 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 84658 0 84714 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 42154 0 42210 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 54390 0 54446 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 65982 0 66038 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 73710 0 73766 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 75642 0 75698 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 77574 0 77630 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 81438 0 81494 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 85302 0 85358 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 87234 0 87290 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 27342 0 27398 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 24766 0 24822 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 360000 400000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 47025570
string GDS_FILE /home/nas163/thkim/efabless/efabless_mpw/openlane/user_proj_example/runs/22_08_29_09_49/results/signoff/user_proj_example.magic.gds
string GDS_START 24451922
<< end >>

