VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO r8_mb8
  CLASS BLOCK ;
  FOREIGN r8_mb8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 132.620 BY 143.340 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END CLK
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 139.340 39.010 143.340 ;
    END
  END RST
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 35.080 10.640 36.680 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 65.440 10.640 67.040 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 95.800 10.640 97.400 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.160 10.640 127.760 130.800 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.900 10.640 21.500 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.260 10.640 51.860 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 80.620 10.640 82.220 130.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.980 10.640 112.580 130.800 ;
    END
  END VPWR
  PIN mx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END mx[0]
  PIN mx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 139.340 119.510 143.340 ;
    END
  END mx[1]
  PIN mx[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 139.340 6.810 143.340 ;
    END
  END mx[2]
  PIN mx[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 139.340 103.410 143.340 ;
    END
  END mx[3]
  PIN mx[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END mx[4]
  PIN mx[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mx[5]
  PIN mx[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 91.840 132.620 92.440 ;
    END
  END mx[6]
  PIN mx[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END mx[7]
  PIN my[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END my[0]
  PIN my[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 108.840 132.620 109.440 ;
    END
  END my[1]
  PIN my[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 74.840 132.620 75.440 ;
    END
  END my[2]
  PIN my[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END my[3]
  PIN my[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 139.340 87.310 143.340 ;
    END
  END my[4]
  PIN my[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 139.340 22.910 143.340 ;
    END
  END my[5]
  PIN my[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END my[6]
  PIN my[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 23.840 132.620 24.440 ;
    END
  END my[7]
  PIN product_final[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END product_final[0]
  PIN product_final[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 139.340 132.390 143.340 ;
    END
  END product_final[10]
  PIN product_final[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 6.840 132.620 7.440 ;
    END
  END product_final[11]
  PIN product_final[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END product_final[12]
  PIN product_final[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END product_final[13]
  PIN product_final[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END product_final[14]
  PIN product_final[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 40.840 132.620 41.440 ;
    END
  END product_final[15]
  PIN product_final[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END product_final[1]
  PIN product_final[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END product_final[2]
  PIN product_final[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 125.840 132.620 126.440 ;
    END
  END product_final[3]
  PIN product_final[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 139.340 55.110 143.340 ;
    END
  END product_final[4]
  PIN product_final[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 139.340 71.210 143.340 ;
    END
  END product_final[5]
  PIN product_final[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END product_final[6]
  PIN product_final[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END product_final[7]
  PIN product_final[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END product_final[8]
  PIN product_final[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 128.620 57.840 132.620 58.440 ;
    END
  END product_final[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 126.960 130.645 ;
      LAYER met1 ;
        RECT 0.070 10.640 132.410 130.800 ;
      LAYER met2 ;
        RECT 0.100 139.060 6.250 139.340 ;
        RECT 7.090 139.060 22.350 139.340 ;
        RECT 23.190 139.060 38.450 139.340 ;
        RECT 39.290 139.060 54.550 139.340 ;
        RECT 55.390 139.060 70.650 139.340 ;
        RECT 71.490 139.060 86.750 139.340 ;
        RECT 87.590 139.060 102.850 139.340 ;
        RECT 103.690 139.060 118.950 139.340 ;
        RECT 119.790 139.060 131.830 139.340 ;
        RECT 0.100 4.280 132.380 139.060 ;
        RECT 0.650 3.670 12.690 4.280 ;
        RECT 13.530 3.670 28.790 4.280 ;
        RECT 29.630 3.670 44.890 4.280 ;
        RECT 45.730 3.670 60.990 4.280 ;
        RECT 61.830 3.670 77.090 4.280 ;
        RECT 77.930 3.670 93.190 4.280 ;
        RECT 94.030 3.670 109.290 4.280 ;
        RECT 110.130 3.670 125.390 4.280 ;
        RECT 126.230 3.670 132.380 4.280 ;
      LAYER met3 ;
        RECT 4.400 132.240 129.410 133.105 ;
        RECT 4.000 126.840 129.410 132.240 ;
        RECT 4.000 125.440 128.220 126.840 ;
        RECT 4.000 116.640 129.410 125.440 ;
        RECT 4.400 115.240 129.410 116.640 ;
        RECT 4.000 109.840 129.410 115.240 ;
        RECT 4.000 108.440 128.220 109.840 ;
        RECT 4.000 99.640 129.410 108.440 ;
        RECT 4.400 98.240 129.410 99.640 ;
        RECT 4.000 92.840 129.410 98.240 ;
        RECT 4.000 91.440 128.220 92.840 ;
        RECT 4.000 82.640 129.410 91.440 ;
        RECT 4.400 81.240 129.410 82.640 ;
        RECT 4.000 75.840 129.410 81.240 ;
        RECT 4.000 74.440 128.220 75.840 ;
        RECT 4.000 65.640 129.410 74.440 ;
        RECT 4.400 64.240 129.410 65.640 ;
        RECT 4.000 58.840 129.410 64.240 ;
        RECT 4.000 57.440 128.220 58.840 ;
        RECT 4.000 48.640 129.410 57.440 ;
        RECT 4.400 47.240 129.410 48.640 ;
        RECT 4.000 41.840 129.410 47.240 ;
        RECT 4.000 40.440 128.220 41.840 ;
        RECT 4.000 31.640 129.410 40.440 ;
        RECT 4.400 30.240 129.410 31.640 ;
        RECT 4.000 24.840 129.410 30.240 ;
        RECT 4.000 23.440 128.220 24.840 ;
        RECT 4.000 14.640 129.410 23.440 ;
        RECT 4.400 13.240 129.410 14.640 ;
        RECT 4.000 7.840 129.410 13.240 ;
        RECT 4.000 6.975 128.220 7.840 ;
  END
END r8_mb8
END LIBRARY

