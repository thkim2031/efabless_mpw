VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sa_2D
  CLASS BLOCK ;
  FOREIGN sa_2D ;
  ORIGIN 0.000 0.000 ;
  SIZE 210.460 BY 221.180 ;
  PIN AA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END AA[0]
  PIN AA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END AA[1]
  PIN AA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END AA[2]
  PIN AA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END AA[3]
  PIN AA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 217.180 16.470 221.180 ;
    END
  END AA[4]
  PIN AA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 81.640 210.460 82.240 ;
    END
  END AA[5]
  PIN AA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 217.180 177.470 221.180 ;
    END
  END AA[6]
  PIN AA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 217.180 0.370 221.180 ;
    END
  END AA[7]
  PIN BB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 13.640 210.460 14.240 ;
    END
  END BB[0]
  PIN BB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 217.180 145.270 221.180 ;
    END
  END BB[1]
  PIN BB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END BB[2]
  PIN BB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END BB[3]
  PIN BB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 30.640 210.460 31.240 ;
    END
  END BB[4]
  PIN BB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 217.180 32.570 221.180 ;
    END
  END BB[5]
  PIN BB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 47.640 210.460 48.240 ;
    END
  END BB[6]
  PIN BB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END BB[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 217.180 96.970 221.180 ;
    END
  END CLK
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END RST
  PIN SHIFTEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END SHIFTEN[0]
  PIN SHIFTEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END SHIFTEN[1]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 209.680 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 209.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 209.680 ;
    END
  END VPWR
  PIN Y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END Y[0]
  PIN Y[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END Y[10]
  PIN Y[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 149.640 210.460 150.240 ;
    END
  END Y[11]
  PIN Y[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END Y[12]
  PIN Y[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 217.180 129.170 221.180 ;
    END
  END Y[13]
  PIN Y[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 217.180 80.870 221.180 ;
    END
  END Y[14]
  PIN Y[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 200.640 210.460 201.240 ;
    END
  END Y[15]
  PIN Y[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 166.640 210.460 167.240 ;
    END
  END Y[16]
  PIN Y[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 115.640 210.460 116.240 ;
    END
  END Y[17]
  PIN Y[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 217.180 161.370 221.180 ;
    END
  END Y[18]
  PIN Y[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END Y[19]
  PIN Y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END Y[1]
  PIN Y[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END Y[20]
  PIN Y[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 183.640 210.460 184.240 ;
    END
  END Y[21]
  PIN Y[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END Y[22]
  PIN Y[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 132.640 210.460 133.240 ;
    END
  END Y[23]
  PIN Y[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END Y[24]
  PIN Y[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 217.180 113.070 221.180 ;
    END
  END Y[25]
  PIN Y[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 64.640 210.460 65.240 ;
    END
  END Y[26]
  PIN Y[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END Y[27]
  PIN Y[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END Y[28]
  PIN Y[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END Y[29]
  PIN Y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END Y[2]
  PIN Y[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END Y[30]
  PIN Y[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 217.180 209.670 221.180 ;
    END
  END Y[31]
  PIN Y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 217.180 193.570 221.180 ;
    END
  END Y[3]
  PIN Y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 217.180 48.670 221.180 ;
    END
  END Y[4]
  PIN Y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 217.180 64.770 221.180 ;
    END
  END Y[5]
  PIN Y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END Y[6]
  PIN Y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END Y[7]
  PIN Y[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END Y[8]
  PIN Y[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 206.460 98.640 210.460 99.240 ;
    END
  END Y[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 204.700 209.525 ;
      LAYER met1 ;
        RECT 0.070 9.560 209.690 209.680 ;
      LAYER met2 ;
        RECT 0.650 216.900 15.910 217.180 ;
        RECT 16.750 216.900 32.010 217.180 ;
        RECT 32.850 216.900 48.110 217.180 ;
        RECT 48.950 216.900 64.210 217.180 ;
        RECT 65.050 216.900 80.310 217.180 ;
        RECT 81.150 216.900 96.410 217.180 ;
        RECT 97.250 216.900 112.510 217.180 ;
        RECT 113.350 216.900 128.610 217.180 ;
        RECT 129.450 216.900 144.710 217.180 ;
        RECT 145.550 216.900 160.810 217.180 ;
        RECT 161.650 216.900 176.910 217.180 ;
        RECT 177.750 216.900 193.010 217.180 ;
        RECT 193.850 216.900 209.110 217.180 ;
        RECT 0.100 4.280 209.660 216.900 ;
        RECT 0.650 4.000 15.910 4.280 ;
        RECT 16.750 4.000 32.010 4.280 ;
        RECT 32.850 4.000 48.110 4.280 ;
        RECT 48.950 4.000 64.210 4.280 ;
        RECT 65.050 4.000 80.310 4.280 ;
        RECT 81.150 4.000 96.410 4.280 ;
        RECT 97.250 4.000 112.510 4.280 ;
        RECT 113.350 4.000 128.610 4.280 ;
        RECT 129.450 4.000 144.710 4.280 ;
        RECT 145.550 4.000 160.810 4.280 ;
        RECT 161.650 4.000 176.910 4.280 ;
        RECT 177.750 4.000 193.010 4.280 ;
        RECT 193.850 4.000 209.110 4.280 ;
      LAYER met3 ;
        RECT 4.000 205.040 206.460 209.605 ;
        RECT 4.400 203.640 206.460 205.040 ;
        RECT 4.000 201.640 206.460 203.640 ;
        RECT 4.000 200.240 206.060 201.640 ;
        RECT 4.000 188.040 206.460 200.240 ;
        RECT 4.400 186.640 206.460 188.040 ;
        RECT 4.000 184.640 206.460 186.640 ;
        RECT 4.000 183.240 206.060 184.640 ;
        RECT 4.000 171.040 206.460 183.240 ;
        RECT 4.400 169.640 206.460 171.040 ;
        RECT 4.000 167.640 206.460 169.640 ;
        RECT 4.000 166.240 206.060 167.640 ;
        RECT 4.000 154.040 206.460 166.240 ;
        RECT 4.400 152.640 206.460 154.040 ;
        RECT 4.000 150.640 206.460 152.640 ;
        RECT 4.000 149.240 206.060 150.640 ;
        RECT 4.000 137.040 206.460 149.240 ;
        RECT 4.400 135.640 206.460 137.040 ;
        RECT 4.000 133.640 206.460 135.640 ;
        RECT 4.000 132.240 206.060 133.640 ;
        RECT 4.000 120.040 206.460 132.240 ;
        RECT 4.400 118.640 206.460 120.040 ;
        RECT 4.000 116.640 206.460 118.640 ;
        RECT 4.000 115.240 206.060 116.640 ;
        RECT 4.000 103.040 206.460 115.240 ;
        RECT 4.400 101.640 206.460 103.040 ;
        RECT 4.000 99.640 206.460 101.640 ;
        RECT 4.000 98.240 206.060 99.640 ;
        RECT 4.000 86.040 206.460 98.240 ;
        RECT 4.400 84.640 206.460 86.040 ;
        RECT 4.000 82.640 206.460 84.640 ;
        RECT 4.000 81.240 206.060 82.640 ;
        RECT 4.000 69.040 206.460 81.240 ;
        RECT 4.400 67.640 206.460 69.040 ;
        RECT 4.000 65.640 206.460 67.640 ;
        RECT 4.000 64.240 206.060 65.640 ;
        RECT 4.000 52.040 206.460 64.240 ;
        RECT 4.400 50.640 206.460 52.040 ;
        RECT 4.000 48.640 206.460 50.640 ;
        RECT 4.000 47.240 206.060 48.640 ;
        RECT 4.000 35.040 206.460 47.240 ;
        RECT 4.400 33.640 206.460 35.040 ;
        RECT 4.000 31.640 206.460 33.640 ;
        RECT 4.000 30.240 206.060 31.640 ;
        RECT 4.000 18.040 206.460 30.240 ;
        RECT 4.400 16.640 206.460 18.040 ;
        RECT 4.000 14.640 206.460 16.640 ;
        RECT 4.000 13.240 206.060 14.640 ;
        RECT 4.000 10.715 206.460 13.240 ;
  END
END sa_2D
END LIBRARY

