
  //######################//
 // 	CLA Parameters      //
//######################//
//for test bench
`define P_W 16
parameter N=16;

//for main module
parameter N_16=16;
parameter WIDTH=32;



