VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLA_16
  CLASS BLOCK ;
  FOREIGN CLA_16 ;
  ORIGIN 0.000 0.000 ;
  SIZE 88.600 BY 99.320 ;
  PIN CIN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END CIN
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END CLK
  PIN COUT_FINAL
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END COUT_FINAL
  PIN OPA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END OPA[0]
  PIN OPA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 95.320 3.590 99.320 ;
    END
  END OPA[10]
  PIN OPA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 40.840 88.600 41.440 ;
    END
  END OPA[11]
  PIN OPA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 95.320 74.430 99.320 ;
    END
  END OPA[12]
  PIN OPA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END OPA[13]
  PIN OPA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 10.240 88.600 10.840 ;
    END
  END OPA[14]
  PIN OPA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 95.320 61.550 99.320 ;
    END
  END OPA[15]
  PIN OPA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 3.440 88.600 4.040 ;
    END
  END OPA[1]
  PIN OPA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END OPA[2]
  PIN OPA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 17.040 88.600 17.640 ;
    END
  END OPA[3]
  PIN OPA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 95.320 10.030 99.320 ;
    END
  END OPA[4]
  PIN OPA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 23.840 88.600 24.440 ;
    END
  END OPA[5]
  PIN OPA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END OPA[6]
  PIN OPA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 95.320 39.010 99.320 ;
    END
  END OPA[7]
  PIN OPA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END OPA[8]
  PIN OPA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END OPA[9]
  PIN OPB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END OPB[0]
  PIN OPB[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END OPB[10]
  PIN OPB[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END OPB[11]
  PIN OPB[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 71.440 88.600 72.040 ;
    END
  END OPB[12]
  PIN OPB[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END OPB[13]
  PIN OPB[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 95.320 51.890 99.320 ;
    END
  END OPB[14]
  PIN OPB[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 95.320 32.570 99.320 ;
    END
  END OPB[15]
  PIN OPB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 91.840 88.600 92.440 ;
    END
  END OPB[1]
  PIN OPB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 78.240 88.600 78.840 ;
    END
  END OPB[2]
  PIN OPB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 54.440 88.600 55.040 ;
    END
  END OPB[3]
  PIN OPB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 95.320 67.990 99.320 ;
    END
  END OPB[4]
  PIN OPB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END OPB[5]
  PIN OPB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END OPB[6]
  PIN OPB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END OPB[7]
  PIN OPB[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 85.040 88.600 85.640 ;
    END
  END OPB[8]
  PIN OPB[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END OPB[9]
  PIN PHI
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 61.240 88.600 61.840 ;
    END
  END PHI
  PIN SUM_FINAL[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END SUM_FINAL[0]
  PIN SUM_FINAL[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 95.320 45.450 99.320 ;
    END
  END SUM_FINAL[10]
  PIN SUM_FINAL[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 30.640 88.600 31.240 ;
    END
  END SUM_FINAL[11]
  PIN SUM_FINAL[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END SUM_FINAL[12]
  PIN SUM_FINAL[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END SUM_FINAL[13]
  PIN SUM_FINAL[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END SUM_FINAL[14]
  PIN SUM_FINAL[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END SUM_FINAL[15]
  PIN SUM_FINAL[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END SUM_FINAL[1]
  PIN SUM_FINAL[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 95.320 87.310 99.320 ;
    END
  END SUM_FINAL[2]
  PIN SUM_FINAL[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 95.320 80.870 99.320 ;
    END
  END SUM_FINAL[3]
  PIN SUM_FINAL[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 95.320 16.470 99.320 ;
    END
  END SUM_FINAL[4]
  PIN SUM_FINAL[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 95.320 22.910 99.320 ;
    END
  END SUM_FINAL[5]
  PIN SUM_FINAL[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END SUM_FINAL[6]
  PIN SUM_FINAL[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END SUM_FINAL[7]
  PIN SUM_FINAL[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END SUM_FINAL[8]
  PIN SUM_FINAL[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 84.600 47.640 88.600 48.240 ;
    END
  END SUM_FINAL[9]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.040 10.640 25.640 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.360 10.640 44.960 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 62.680 10.640 64.280 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.000 10.640 83.600 87.280 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 14.380 10.640 15.980 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.700 10.640 35.300 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.020 10.640 54.620 87.280 ;
    END
    PORT
      LAYER met4 ;
        RECT 72.340 10.640 73.940 87.280 ;
    END
  END VPWR
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 82.800 87.125 ;
      LAYER met1 ;
        RECT 0.070 10.240 87.330 87.280 ;
      LAYER met2 ;
        RECT 0.100 95.040 3.030 95.725 ;
        RECT 3.870 95.040 9.470 95.725 ;
        RECT 10.310 95.040 15.910 95.725 ;
        RECT 16.750 95.040 22.350 95.725 ;
        RECT 23.190 95.040 32.010 95.725 ;
        RECT 32.850 95.040 38.450 95.725 ;
        RECT 39.290 95.040 44.890 95.725 ;
        RECT 45.730 95.040 51.330 95.725 ;
        RECT 52.170 95.040 60.990 95.725 ;
        RECT 61.830 95.040 67.430 95.725 ;
        RECT 68.270 95.040 73.870 95.725 ;
        RECT 74.710 95.040 80.310 95.725 ;
        RECT 81.150 95.040 86.750 95.725 ;
        RECT 0.100 4.280 87.300 95.040 ;
        RECT 0.650 3.555 6.250 4.280 ;
        RECT 7.090 3.555 12.690 4.280 ;
        RECT 13.530 3.555 19.130 4.280 ;
        RECT 19.970 3.555 25.570 4.280 ;
        RECT 26.410 3.555 35.230 4.280 ;
        RECT 36.070 3.555 41.670 4.280 ;
        RECT 42.510 3.555 48.110 4.280 ;
        RECT 48.950 3.555 54.550 4.280 ;
        RECT 55.390 3.555 64.210 4.280 ;
        RECT 65.050 3.555 70.650 4.280 ;
        RECT 71.490 3.555 77.090 4.280 ;
        RECT 77.930 3.555 83.530 4.280 ;
        RECT 84.370 3.555 87.300 4.280 ;
      LAYER met3 ;
        RECT 4.400 94.840 85.250 95.705 ;
        RECT 4.000 92.840 85.250 94.840 ;
        RECT 4.000 91.440 84.200 92.840 ;
        RECT 4.000 89.440 85.250 91.440 ;
        RECT 4.400 88.040 85.250 89.440 ;
        RECT 4.000 86.040 85.250 88.040 ;
        RECT 4.000 84.640 84.200 86.040 ;
        RECT 4.000 82.640 85.250 84.640 ;
        RECT 4.400 81.240 85.250 82.640 ;
        RECT 4.000 79.240 85.250 81.240 ;
        RECT 4.000 77.840 84.200 79.240 ;
        RECT 4.000 75.840 85.250 77.840 ;
        RECT 4.400 74.440 85.250 75.840 ;
        RECT 4.000 72.440 85.250 74.440 ;
        RECT 4.000 71.040 84.200 72.440 ;
        RECT 4.000 69.040 85.250 71.040 ;
        RECT 4.400 67.640 85.250 69.040 ;
        RECT 4.000 62.240 85.250 67.640 ;
        RECT 4.000 60.840 84.200 62.240 ;
        RECT 4.000 58.840 85.250 60.840 ;
        RECT 4.400 57.440 85.250 58.840 ;
        RECT 4.000 55.440 85.250 57.440 ;
        RECT 4.000 54.040 84.200 55.440 ;
        RECT 4.000 52.040 85.250 54.040 ;
        RECT 4.400 50.640 85.250 52.040 ;
        RECT 4.000 48.640 85.250 50.640 ;
        RECT 4.000 47.240 84.200 48.640 ;
        RECT 4.000 45.240 85.250 47.240 ;
        RECT 4.400 43.840 85.250 45.240 ;
        RECT 4.000 41.840 85.250 43.840 ;
        RECT 4.000 40.440 84.200 41.840 ;
        RECT 4.000 38.440 85.250 40.440 ;
        RECT 4.400 37.040 85.250 38.440 ;
        RECT 4.000 31.640 85.250 37.040 ;
        RECT 4.000 30.240 84.200 31.640 ;
        RECT 4.000 28.240 85.250 30.240 ;
        RECT 4.400 26.840 85.250 28.240 ;
        RECT 4.000 24.840 85.250 26.840 ;
        RECT 4.000 23.440 84.200 24.840 ;
        RECT 4.000 21.440 85.250 23.440 ;
        RECT 4.400 20.040 85.250 21.440 ;
        RECT 4.000 18.040 85.250 20.040 ;
        RECT 4.000 16.640 84.200 18.040 ;
        RECT 4.000 14.640 85.250 16.640 ;
        RECT 4.400 13.240 85.250 14.640 ;
        RECT 4.000 11.240 85.250 13.240 ;
        RECT 4.000 9.840 84.200 11.240 ;
        RECT 4.000 7.840 85.250 9.840 ;
        RECT 4.400 6.440 85.250 7.840 ;
        RECT 4.000 4.440 85.250 6.440 ;
        RECT 4.000 3.575 84.200 4.440 ;
  END
END CLA_16
END LIBRARY

