VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sa_2D
  CLASS BLOCK ;
  FOREIGN sa_2D ;
  ORIGIN 0.000 0.000 ;
  SIZE 187.305 BY 198.025 ;
  PIN AA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END AA[0]
  PIN AA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END AA[1]
  PIN AA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END AA[2]
  PIN AA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END AA[3]
  PIN AA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 194.025 13.250 198.025 ;
    END
  END AA[4]
  PIN AA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 74.840 187.305 75.440 ;
    END
  END AA[5]
  PIN AA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 194.025 158.150 198.025 ;
    END
  END AA[6]
  PIN AA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END AA[7]
  PIN BB[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 13.640 187.305 14.240 ;
    END
  END BB[0]
  PIN BB[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 194.025 129.170 198.025 ;
    END
  END BB[1]
  PIN BB[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 0.040 187.305 0.640 ;
    END
  END BB[2]
  PIN BB[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END BB[3]
  PIN BB[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 30.640 187.305 31.240 ;
    END
  END BB[4]
  PIN BB[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 194.025 29.350 198.025 ;
    END
  END BB[5]
  PIN BB[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 44.240 187.305 44.840 ;
    END
  END BB[6]
  PIN BB[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END BB[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 194.025 87.310 198.025 ;
    END
  END CLK
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END RST
  PIN SHIFTEN[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END SHIFTEN[0]
  PIN SHIFTEN[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END SHIFTEN[1]
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 185.200 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 185.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 185.200 ;
    END
  END VPWR
  PIN Y[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END Y[0]
  PIN Y[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END Y[10]
  PIN Y[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 136.040 187.305 136.640 ;
    END
  END Y[11]
  PIN Y[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END Y[12]
  PIN Y[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 194.025 116.290 198.025 ;
    END
  END Y[13]
  PIN Y[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 194.025 71.210 198.025 ;
    END
  END Y[14]
  PIN Y[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 183.640 187.305 184.240 ;
    END
  END Y[15]
  PIN Y[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 153.040 187.305 153.640 ;
    END
  END Y[16]
  PIN Y[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 105.440 187.305 106.040 ;
    END
  END Y[17]
  PIN Y[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 194.025 145.270 198.025 ;
    END
  END Y[18]
  PIN Y[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END Y[19]
  PIN Y[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END Y[1]
  PIN Y[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END Y[20]
  PIN Y[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 166.640 187.305 167.240 ;
    END
  END Y[21]
  PIN Y[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END Y[22]
  PIN Y[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 122.440 187.305 123.040 ;
    END
  END Y[23]
  PIN Y[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END Y[24]
  PIN Y[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 194.025 100.190 198.025 ;
    END
  END Y[25]
  PIN Y[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 61.240 187.305 61.840 ;
    END
  END Y[26]
  PIN Y[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END Y[27]
  PIN Y[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END Y[28]
  PIN Y[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END Y[29]
  PIN Y[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END Y[2]
  PIN Y[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END Y[30]
  PIN Y[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 194.025 187.130 198.025 ;
    END
  END Y[31]
  PIN Y[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 194.025 174.250 198.025 ;
    END
  END Y[3]
  PIN Y[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 194.025 42.230 198.025 ;
    END
  END Y[4]
  PIN Y[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 194.025 58.330 198.025 ;
    END
  END Y[5]
  PIN Y[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END Y[6]
  PIN Y[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END Y[7]
  PIN Y[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END Y[8]
  PIN Y[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 183.305 91.840 187.305 92.440 ;
    END
  END Y[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 181.700 185.045 ;
      LAYER met1 ;
        RECT 0.070 9.560 187.150 185.200 ;
      LAYER met2 ;
        RECT 0.100 193.745 12.690 197.725 ;
        RECT 13.530 193.745 28.790 197.725 ;
        RECT 29.630 193.745 41.670 197.725 ;
        RECT 42.510 193.745 57.770 197.725 ;
        RECT 58.610 193.745 70.650 197.725 ;
        RECT 71.490 193.745 86.750 197.725 ;
        RECT 87.590 193.745 99.630 197.725 ;
        RECT 100.470 193.745 115.730 197.725 ;
        RECT 116.570 193.745 128.610 197.725 ;
        RECT 129.450 193.745 144.710 197.725 ;
        RECT 145.550 193.745 157.590 197.725 ;
        RECT 158.430 193.745 173.690 197.725 ;
        RECT 174.530 193.745 186.570 197.725 ;
        RECT 0.100 4.280 187.120 193.745 ;
        RECT 0.650 0.155 12.690 4.280 ;
        RECT 13.530 0.155 28.790 4.280 ;
        RECT 29.630 0.155 41.670 4.280 ;
        RECT 42.510 0.155 57.770 4.280 ;
        RECT 58.610 0.155 70.650 4.280 ;
        RECT 71.490 0.155 86.750 4.280 ;
        RECT 87.590 0.155 99.630 4.280 ;
        RECT 100.470 0.155 115.730 4.280 ;
        RECT 116.570 0.155 128.610 4.280 ;
        RECT 129.450 0.155 144.710 4.280 ;
        RECT 145.550 0.155 157.590 4.280 ;
        RECT 158.430 0.155 173.690 4.280 ;
        RECT 174.530 0.155 187.120 4.280 ;
      LAYER met3 ;
        RECT 4.400 196.840 183.305 197.705 ;
        RECT 4.000 184.640 183.305 196.840 ;
        RECT 4.400 183.240 182.905 184.640 ;
        RECT 4.000 167.640 183.305 183.240 ;
        RECT 4.400 166.240 182.905 167.640 ;
        RECT 4.000 154.040 183.305 166.240 ;
        RECT 4.400 152.640 182.905 154.040 ;
        RECT 4.000 137.040 183.305 152.640 ;
        RECT 4.400 135.640 182.905 137.040 ;
        RECT 4.000 123.440 183.305 135.640 ;
        RECT 4.400 122.040 182.905 123.440 ;
        RECT 4.000 106.440 183.305 122.040 ;
        RECT 4.400 105.040 182.905 106.440 ;
        RECT 4.000 92.840 183.305 105.040 ;
        RECT 4.400 91.440 182.905 92.840 ;
        RECT 4.000 75.840 183.305 91.440 ;
        RECT 4.400 74.440 182.905 75.840 ;
        RECT 4.000 62.240 183.305 74.440 ;
        RECT 4.400 60.840 182.905 62.240 ;
        RECT 4.000 45.240 183.305 60.840 ;
        RECT 4.400 43.840 182.905 45.240 ;
        RECT 4.000 31.640 183.305 43.840 ;
        RECT 4.400 30.240 182.905 31.640 ;
        RECT 4.000 14.640 183.305 30.240 ;
        RECT 4.400 13.240 182.905 14.640 ;
        RECT 4.000 1.040 183.305 13.240 ;
        RECT 4.000 0.175 182.905 1.040 ;
      LAYER met4 ;
        RECT 87.695 15.135 88.025 160.305 ;
  END
END sa_2D
END LIBRARY

