VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO r8_mb8
  CLASS BLOCK ;
  FOREIGN r8_mb8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 122.630 BY 133.350 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END CLK
  PIN RST
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 129.350 32.570 133.350 ;
    END
  END RST
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 32.550 10.640 34.150 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 60.380 10.640 61.980 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.210 10.640 89.810 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 116.040 10.640 117.640 122.640 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.635 10.640 20.235 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.465 10.640 48.065 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.295 10.640 75.895 122.640 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.125 10.640 103.725 122.640 ;
    END
  END VPWR
  PIN mx[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END mx[0]
  PIN mx[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 129.350 106.630 133.350 ;
    END
  END mx[1]
  PIN mx[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 129.350 3.590 133.350 ;
    END
  END mx[2]
  PIN mx[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 129.350 90.530 133.350 ;
    END
  END mx[3]
  PIN mx[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END mx[4]
  PIN mx[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mx[5]
  PIN mx[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 88.440 122.630 89.040 ;
    END
  END mx[6]
  PIN mx[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END mx[7]
  PIN my[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END my[0]
  PIN my[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 102.040 122.630 102.640 ;
    END
  END my[1]
  PIN my[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 71.440 122.630 72.040 ;
    END
  END my[2]
  PIN my[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END my[3]
  PIN my[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 129.350 77.650 133.350 ;
    END
  END my[4]
  PIN my[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 129.350 16.470 133.350 ;
    END
  END my[5]
  PIN my[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END my[6]
  PIN my[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 23.840 122.630 24.440 ;
    END
  END my[7]
  PIN product_final[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END product_final[0]
  PIN product_final[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 129.350 119.510 133.350 ;
    END
  END product_final[10]
  PIN product_final[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 10.240 122.630 10.840 ;
    END
  END product_final[11]
  PIN product_final[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END product_final[12]
  PIN product_final[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END product_final[13]
  PIN product_final[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END product_final[14]
  PIN product_final[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 40.840 122.630 41.440 ;
    END
  END product_final[15]
  PIN product_final[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END product_final[1]
  PIN product_final[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END product_final[2]
  PIN product_final[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 119.040 122.630 119.640 ;
    END
  END product_final[3]
  PIN product_final[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 129.350 48.670 133.350 ;
    END
  END product_final[4]
  PIN product_final[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 129.350 61.550 133.350 ;
    END
  END product_final[5]
  PIN product_final[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END product_final[6]
  PIN product_final[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END product_final[7]
  PIN product_final[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END product_final[8]
  PIN product_final[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 118.630 57.840 122.630 58.440 ;
    END
  END product_final[9]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 116.840 122.485 ;
      LAYER met1 ;
        RECT 0.070 10.640 119.530 122.640 ;
      LAYER met2 ;
        RECT 0.100 129.070 3.030 129.350 ;
        RECT 3.870 129.070 15.910 129.350 ;
        RECT 16.750 129.070 32.010 129.350 ;
        RECT 32.850 129.070 48.110 129.350 ;
        RECT 48.950 129.070 60.990 129.350 ;
        RECT 61.830 129.070 77.090 129.350 ;
        RECT 77.930 129.070 89.970 129.350 ;
        RECT 90.810 129.070 106.070 129.350 ;
        RECT 106.910 129.070 118.950 129.350 ;
        RECT 0.100 4.280 119.500 129.070 ;
        RECT 0.650 4.000 12.690 4.280 ;
        RECT 13.530 4.000 28.790 4.280 ;
        RECT 29.630 4.000 41.670 4.280 ;
        RECT 42.510 4.000 57.770 4.280 ;
        RECT 58.610 4.000 70.650 4.280 ;
        RECT 71.490 4.000 86.750 4.280 ;
        RECT 87.590 4.000 102.850 4.280 ;
        RECT 103.690 4.000 115.730 4.280 ;
        RECT 116.570 4.000 119.500 4.280 ;
      LAYER met3 ;
        RECT 4.400 122.040 119.290 122.905 ;
        RECT 4.000 120.040 119.290 122.040 ;
        RECT 4.000 118.640 118.230 120.040 ;
        RECT 4.000 109.840 119.290 118.640 ;
        RECT 4.400 108.440 119.290 109.840 ;
        RECT 4.000 103.040 119.290 108.440 ;
        RECT 4.000 101.640 118.230 103.040 ;
        RECT 4.000 92.840 119.290 101.640 ;
        RECT 4.400 91.440 119.290 92.840 ;
        RECT 4.000 89.440 119.290 91.440 ;
        RECT 4.000 88.040 118.230 89.440 ;
        RECT 4.000 75.840 119.290 88.040 ;
        RECT 4.400 74.440 119.290 75.840 ;
        RECT 4.000 72.440 119.290 74.440 ;
        RECT 4.000 71.040 118.230 72.440 ;
        RECT 4.000 62.240 119.290 71.040 ;
        RECT 4.400 60.840 119.290 62.240 ;
        RECT 4.000 58.840 119.290 60.840 ;
        RECT 4.000 57.440 118.230 58.840 ;
        RECT 4.000 45.240 119.290 57.440 ;
        RECT 4.400 43.840 119.290 45.240 ;
        RECT 4.000 41.840 119.290 43.840 ;
        RECT 4.000 40.440 118.230 41.840 ;
        RECT 4.000 31.640 119.290 40.440 ;
        RECT 4.400 30.240 119.290 31.640 ;
        RECT 4.000 24.840 119.290 30.240 ;
        RECT 4.000 23.440 118.230 24.840 ;
        RECT 4.000 14.640 119.290 23.440 ;
        RECT 4.400 13.240 119.290 14.640 ;
        RECT 4.000 11.240 119.290 13.240 ;
        RECT 4.000 10.715 118.230 11.240 ;
  END
END r8_mb8
END LIBRARY

